package riscv_test_pkg;

  import opcodes::*;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "exec_record.svh"
  `include "opcode_seq_item.svh"
  `include "iss_class.svh"

  `include "riscv_monitor.svh"
  `include "riscv_tracer.svh"
  `include "riscv_scoreboard.svh"
  `include "riscv_coverage.svh"

  `include "execute_driver.svh"
  `include "execute_agent.svh"
  `include "execute_env.svh"
  `include "execute_test.svh"

  // tests derived from execute_test

  `include "mem_test.svh"
  `include "fibonacci.svh"
  
endpackage
